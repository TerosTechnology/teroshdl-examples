module evaluate_example();

// Unsigned binary: 3
localparam [2:0] e_binary_unsigned = 3'b011;
// Signed binary 7 (unsigned), -1 (signed)
localparam [2:0] e_binary_signed = 3'b111;
// Unsigned octal 19
localparam [5:0] e_octal = 6'o23;
// Unsigned hexadecimal 35
localparam [5:0] e_hex = 6'h23                                              ;

endmodule

